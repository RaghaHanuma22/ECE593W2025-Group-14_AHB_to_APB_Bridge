// File: ahb_apb_assertions.sv
`include "uvm_macros.svh"
import uvm_pkg::*;

module ahb_apb_assertions (
    // AHB and APB interfaces
    input logic Hclk, Hresetn, Hwrite, Hreadyin, Hreadyout,
    input logic [1:0] Htrans, input logic [31:0] Hwdata, Haddr,
    input logic [1:0] Hresp, input logic Pwrite, input logic [2:0] Pselx,
    input logic Penable, input logic [31:0] Paddr, Pwdata, Prdata,
    input logic valid, input logic [31:0] Haddr1, Haddr2, input logic Hwritereg
);

    //////////////////////////////////////////////////////////////////
    // 1. AHB Protocol Assertions
    //////////////////////////////////////////////////////////////////
    
    // Valid HTRANS values check
    property valid_htrans_p;
        @(posedge Hclk) disable iff (!Hresetn)
        $isunknown(Htrans) == 0 |-> Htrans inside {2'b00, 2'b10, 2'b11};
    endproperty
    
    VALID_HTRANS: assert property(valid_htrans_p)
        else `uvm_error("VALID_HTRANS", $sformatf("Invalid HTRANS value detected: %b at time %0t", Htrans, $time))
    
    cover property(@(posedge Hclk) (Htrans == 2'b00))
        $info("HTRANS IDLE covered");
    cover property(@(posedge Hclk) (Htrans == 2'b10))
        $info("HTRANS NONSEQ covered");
    
    // Hresp should be OKAY during normal operation
    property hresp_okay_p;
        @(posedge Hclk) disable iff (!Hresetn)
        1'b1 |-> Hresp == 2'b00;
    endproperty
    
    HRESP_OKAY: assert property(hresp_okay_p)
        else `uvm_error("HRESP_OKAY", $sformatf("HRESP not OKAY during normal operation at time %0t", $time))
    
    cover property(@(posedge Hclk) Hresp == 2'b00)
        $info("HRESP OKAY covered");
    

    //////////////////////////////////////////////////////////////////
    // 4. Data Transfer Assertions 
    //////////////////////////////////////////////////////////////////
    
    // Pipelining check - simplified to just check address pipelining
    property addr_pipelining_p;
        @(posedge Hclk) disable iff (!Hresetn)
         ($past(Hresetn) && Hresetn && $past($isunknown(Haddr)) == 0) |-> (Haddr1 == $past(Haddr));
    endproperty
    
    ADDR_PIPELINING: assert property(addr_pipelining_p)
        else `uvm_error("ADDR_PIPELINING", $sformatf("Address pipelining violation at time %0t", $time))
    
    cover property(@(posedge Hclk) (Haddr1 == $past(Haddr)))
        $info("Address pipelining covered");
    
    // Valid signal generation check (simplified)
    property valid_signal_gen_p;
        @(posedge Hclk) disable iff (!Hresetn)
        (Hreadyin && (Haddr >= 32'h0 && Haddr <= 32'h7ff) && 
         (Htrans == 2'b10 || Htrans == 2'b11)) |-> !valid;
    endproperty
    
    VALID_SIGNAL_GEN: assert property(valid_signal_gen_p)
        else `uvm_error("VALID_SIGNAL_GEN", $sformatf("Valid signal not generated correctly at time %0t", $time))
    
    cover property(@(posedge Hclk) valid)
        $info("Valid signal generation covered");
    
    //////////////////////////////////////////////////////////////////
    // 5. Reset Behavior Assertions 
    //////////////////////////////////////////////////////////////////
    
    // Reset behavior - check specific outputs
    property reset_behavior_p;
        @(posedge Hclk)
        !Hresetn |=> !Penable;
    endproperty
    
    RESET_BEHAVIOR: assert property(reset_behavior_p)
        else `uvm_error("RESET_BEHAVIOR", $sformatf("Incorrect reset behavior at time %0t", $time))
    
    cover property(@(posedge Hclk) !Hresetn ##1 Hresetn)
        $info("Reset sequence covered");
    
    //////////////////////////////////////////////////////////////////
    // 6. Simple Transaction Assertions (Basic transactions)
    //////////////////////////////////////////////////////////////////
    
    // Basic successful write transaction (very simplified sequence)
    property basic_write_p;
        @(posedge Hclk) disable iff (!Hresetn)
        (Hwrite && Htrans == 2'b10) |=> (Htrans == 2'b00) |-> ##[1:10] Hreadyout;
    endproperty
    
    BASIC_WRITE: assert property(basic_write_p)
        else `uvm_error("BASIC_WRITE", $sformatf("Basic write transaction failed at time %0t", $time))
    
    cover property(@(posedge Hclk) (Hwrite && Htrans == 2'b10) ##1 (Htrans == 2'b00) ##[1:10] Hreadyout)
        $info("Basic write transaction covered");
    
    // Basic successful read transaction (very simplified sequence)
    property basic_read_p;
        @(posedge Hclk) disable iff (!Hresetn)
        (!Hwrite && Htrans == 2'b10) |=> (Htrans == 2'b00) |-> ##[1:10] Hreadyout;
    endproperty
    
    BASIC_READ: assert property(basic_read_p)
        else `uvm_error("BASIC_READ", $sformatf("Basic read transaction failed at time %0t", $time))
    
    cover property(@(posedge Hclk) (!Hwrite && Htrans == 2'b10) ##1 (Htrans == 2'b00) ##[1:10] Hreadyout)
        $info("Basic read transaction covered");

endmodule
